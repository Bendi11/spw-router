module OSERDESE2
#(

)
(

);

endmodule;
