module ISERDESE2
#(
    parameter INTERFACE_TYPE="NETWORKING",
    parameter DATA_WIDTH=8
)
(
    input wire RST,
    input wire CLK,
    input wire D,
    output wire Q1,
    output wire Q2,
    output wire Q3,
    output wire Q4,
    output wire Q5,
    output wire Q6,
    output wire Q7,
    output wire Q8
);

endmodule
