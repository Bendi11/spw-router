module OSERDESE2
#(
    parameter DATA_RATE_OQ="SDR",
    parameter DATA_WIDTH=8
)
(
    input wire CLK,
    output wire OQ,
    input wire D1,
    input wire D2,
    input wire D3,
    input wire D4,
    input wire D5,
    input wire D6,
    input wire D7,
    input wire D8
);

endmodule
