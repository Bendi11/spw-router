module OBUFDS(input wire I, output wire O, output wire OB);

endmodule
